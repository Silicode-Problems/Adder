module adder(a, b, sum);

// Your code here

endmodule : adder